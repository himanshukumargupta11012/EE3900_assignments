question 2.8

V1 v1 0 2
V2 v2 0 1
R1 v1 v3 2
R2 v2 v3 1
C1 v3 0 1u ic=0

.tran 100u 5u uic

.control 
run
wrdata 2.8.dat V(v3)
.endc
.end
